// Bluespec types for supporting the RISC-V Formal Interface (RVFI) defined by
// Claire Wolf.
//
// An RVFI port on a micro is also _really useful_ for tests and trace, in
// addition to formal verification.
package Rvfi;

typedef enum {
    UMode = 0,
    SMode = 1,
    MMode = 2
} Priv deriving (Eq, Bits, FShow);

// The single-instruction-retired RVFI output interface expected in Verilog.
(* always_ready, always_enabled *)
interface Rvfi#(numeric type xlen, numeric type ilen);
    method Bool valid;
    method UInt#(64) order;
    method Bit#(ilen) insn;
    method Bool trap;
    method Bool halt;
    method Bool intr;
    method Priv mode;
    method Bit#(2) ixl;

    interface RvfiRegRead#(xlen) rs1;
    interface RvfiRegRead#(xlen) rs2;
    interface RvfiRegWrite#(xlen) rd;

    method Bit#(xlen) pc_rdata;
    method Bit#(xlen) pc_wdata;

    method Bit#(xlen) mem_addr;
    method Bit#(TDiv#(xlen, 8)) mem_rmask;
    method Bit#(TDiv#(xlen, 8)) mem_wmask;
    method Bit#(xlen) mem_rdata;
    method Bit#(xlen) mem_wdata;
endinterface

// Repeated prefixed signals broken out
(* always_ready, always_enabled *)
interface RvfiRegRead#(numeric type xlen);
    method Bit#(5) addr;
    method Bit#(xlen) data;
endinterface

(* always_ready, always_enabled *)
interface RvfiRegWrite#(numeric type xlen);
    method Bit#(5) addr;
    method Bit#(xlen) wdata;
endinterface

// "Emitter" side interface and utility module for convenience.
interface RvfiEmit#(numeric type xlen, numeric type ilen);
    (* always_ready *)
    method Action retire(RvfiRetire#(xlen, ilen) record);
endinterface

function RvfiEmit#(xlen, ilen) noRvfi;
    return (interface RvfiEmit;
        method Action retire(record) = noAction;
    endinterface);
endfunction

interface RvfiPipe#(numeric type xlen, numeric type ilen);
    interface RvfiEmit#(xlen, ilen) in;
    interface Rvfi#(xlen, ilen) out;
endinterface

module mkRvfiPipe (RvfiPipe#(xlen, ilen));
    let record_wire <- mkRWire;
    let retire_counter <- mkReg(0);
    let {urec, uctr} = fromMaybe(?, record_wire.wget);

    interface RvfiEmit in;
        method Action retire(record);
            record_wire.wset(tuple2(record, retire_counter));
            retire_counter <= retire_counter + 1;
        endmethod
    endinterface

    interface Rvfi out;
        method valid = isValid(record_wire.wget);
        method order = uctr;
        method insn = urec.insn;
        method trap = urec.trap;
        method halt = urec.halt;
        method intr = urec.intr;
        method mode = urec.mode;
        method ixl = urec.ixl;

        method pc_rdata = urec.pc_before;
        method pc_wdata = urec.pc_after;

        method mem_addr = urec.mem_addr;
        method mem_rmask = urec.mem_rmask;
        method mem_wmask = urec.mem_wmask;
        method mem_rdata = urec.mem_rdata;
        method mem_wdata = urec.mem_wdata;

        interface RvfiRegRead rs1;
            method addr = tpl_1(urec.rs1);
            method data = tpl_2(urec.rs1);
        endinterface
        interface RvfiRegRead rs2;
            method addr = tpl_1(urec.rs2);
            method data = tpl_2(urec.rs2);
        endinterface
        interface RvfiRegWrite rd;
            method addr = tpl_1(urec.rd);
            method wdata = tpl_2(urec.rd);
        endinterface

    endinterface
endmodule

// Information about retired instruction, packaged as a struct for convenience.
//
// Two signals are missing here:
// - valid is implicit by this struct existing
// - order is generated by a counter in the pipe module and is not a property
//   of the struct itself.
typedef struct {
    Bit#(ilen) insn;
    Bool trap;
    Bool halt;
    Bool intr;
    Priv mode;
    Bit#(2) ixl;

    Tuple2#(Bit#(5), Bit#(xlen)) rs1;
    Tuple2#(Bit#(5), Bit#(xlen)) rs2;
    Tuple2#(Bit#(5), Bit#(xlen)) rd;

    Bit#(xlen) pc_before;
    Bit#(xlen) pc_after;

    Bit#(xlen) mem_addr;
    Bit#(TDiv#(xlen, 8)) mem_rmask;
    Bit#(TDiv#(xlen, 8)) mem_wmask;
    Bit#(xlen) mem_rdata;
    Bit#(xlen) mem_wdata;
} RvfiRetire#(numeric type xlen, numeric type ilen)
deriving (Bits, FShow);

endpackage
